`ifndef memory_mux_include
`define memory_mux_include
// Memory mux Options
`define  MUX_TRAVERSAL   3'b000
`define  MUX_EXECUTE     3'b001
`define  MUX_CELL        3'b010
`define  MUX_INCR        3'b011
`define  MUX_EQUAL       3'b100
`define  MUX_EDITL       3'b101

`endif
