`ifndef traversal_include
`define traversal_include


`endif
